`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO 
// Engineer:  dariomtz
//////////////////////////////////////////////////////////////////////////////////
module display(
    input [3:0] n,
	output [7:0] d
    );

    assign d = (n == 0) 7'b00000000 :
                (n == 8) 7'b11111110;
                      
endmodule