`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO 
// Engineer:  dariomtz
//////////////////////////////////////////////////////////////////////////////////
module top(
    input [7:0] num,
    output [7:0] leds
    );

    assign leds = num;
                                                
endmodule